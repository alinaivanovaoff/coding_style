//-----------------------------------------------------------------------------
// Original Author: Alina Ivanova
// e-mail: alina.al.ivanova@gmail.com
// web: www.alinaivanovaoff.com
// functions_pkg.sv
// Created: 10.26.2016
//
// Functions package.
//
//-----------------------------------------------------------------------------
// Copyright (c) 2016 by Alina Ivanova
//
// This program is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <http://www.gnu.org/licenses/>.
//-----------------------------------------------------------------------------
package functions_pkg;
   function integer clog2(input integer value);
      value -= 1;
      for (clog2 = 0; value > 0; clog2++) begin
         value = value >> 1;
      end
   endfunction: clog2
endpackage: functions_pkg